`include "../include/tune.v"

// Pentevo project (c) NedoPC 2011
//
// atm palette

module video_palette(
);

endmodule

